* 
* No part of this file can be released without the consent of SMIC.
*
* Note: SMIC recommends that users set VNTOL=1E-9 at .option for more smooth convergence.
******************************************************************************************
* 0.18um Mixed Signal 1P6M with MIM Salicide 1.8V/3.3V RF SPICE Model (for HSPICE only)  *
******************************************************************************************
*
* Release version    : 1.9
*
* Release date       : 12/03/2008(dd/mm/yy)
*
* Simulation tool    : Synopsys Star-HSPICE version 2005.9
*
* Model type         :
*   MOSFET           : HSPICE Level 49(BSIM3V3.2)
*   Junction Diode   : HSPICE Level 3
* 
* Model and subcircuit name         :
*   MOSFET           :
*        *------------------------------------------*
*        |     MOSFET model   |   1.8V   |   3.3V   |
*        |==========================================|
*        |        NMOS        |  n18_rf  |  n33_rf  |
*        *------------------------------------------*
*        |       DNWMOS       | dnw18_rf | dnw33_rf |
*        *------------------------------------------*
*        |        PMOS        |  p18_rf  |  p33_rf  |
*        *------------------------------------------*
*
*        *--------------------------------------------------*
*        |     MOSFET subckt  |     1.8V     |    3.3V      |
*        |==================================================|
*        |        NMOS        |  n18_ckt_rf  |  n33_ckt_rf  |
*        *--------------------------------------------------*
*        |       DNWMOS       | dnw18_ckt_rf | dnw33_ckt_rf |
*        *--------------------------------------------------*
*        |        PMOS        |  p18_ckt_rf  |  p33_ckt_rf  |
*        *--------------------------------------------------*
*
*************************
* 1.8V RF NMOS Subcircuit
*************************
* 11=drain, 2=gate, 31=source, 4=bulk
* lr=gate length, wr=finger width, nf=finger number
.subckt n18_ckt_rf 1 2 3 4 lr=l wr=w nf=finger 
*sar=sa sbr=sb sdr=sd
* scalable unit parameter
* euqivalent circuit saclable parameter
.param
+Rg_rf        = 'max(((724.84*pwr(lr*1e6,2)-356.18*lr*1e6+50.477)+(-72.591*pwr(lr*1e6,2)+34.823*lr*1e6-4.3737)*wr*1e6+(-709.9*pwr(lr*1e6,2)+340.42*lr*1e6-49.734)/(wr*1e6))+((-5161.5*pwr(lr*1e6,2)+1999.2*lr*1e6-33.119)+(531.35*pwr(lr*1e6,2)-224.13*lr*1e6+12.828)*wr*1e6+(3902.6*pwr(lr*1e6,2)-164.08*lr*1e6+386.39)/(wr*1e6))/nf,1e-3)'
+Cgd_rf       = 'max((((0.6677*pwr(lr*1e6,2)-0.4222*lr*1e6+0.0529)*pwr(wr*1e6,2)+(-5.7464*pwr(lr*1e6,2)+3.8016*lr*1e6-0.1298)*wr*1e6+(3.275*pwr(lr*1e6,2)-2.272*lr*1e6+0.6075))*nf+((-3.5823*pwr(lr*1e6,2)+2.4353*lr*1e6-0.3546)*pwr(wr*1e6,2)+(30.068*pwr(lr*1e6,2)-20.101*lr*1e6+2.8423)*wr*1e6+(-23.613*pwr(lr*1e6,2)+15.794*lr*1e6-1.9974)))*1e-15, 1e-18)'
+Cgs_rf       = 'max((((0.0651*pwr(lr*1e6,2)-0.0346*lr*1e6+0.004)*pwr(wr*1e6,2)+(-0.701*pwr(lr*1e6,2)+0.3523*lr*1e6-0.0371)*wr*1e6+(1.0807*pwr(lr*1e6,2)-0.5396*lr*1e6+0.061))*pwr(nf,2)+((-0.1448*pwr(lr*1e6,2)-0.1172*lr*1e6+0.0525)*pwr(wr*1e6,2)+(1.1016*pwr(lr*1e6,2)+2.1538*lr*1e6-0.8227)*wr*1e6+(-11.232*pwr(lr*1e6,2)+1.8929*lr*1e6+0.7917))*nf+((-2.1156*pwr(lr*1e6,2)+2.368*lr*1e6-0.5178)*pwr(wr*1e6,2)+(33.552*pwr(lr*1e6,2)-34.449*lr*1e6+6.9433)*wr*1e6+(-54.224*pwr(lr*1e6,2)+52.226*lr*1e6-7.2535)))*1e-15, 1e-18)'
+Cds_rf       = 'max((((1.2656*pwr(lr*1e6,2)-0.8625*lr*1e6+0.1269)*pwr(wr*1e6,2)+(-14.055*pwr(lr*1e6,2)+8.8032*lr*1e6-0.7362)*wr*1e6+(16.189*pwr(lr*1e6,2)-11.156*lr*1e6+1.6503))*nf+((-6.6026*pwr(lr*1e6,2)+3.9526*lr*1e6-0.3798)*pwr(wr*1e6,2)+(76.57*pwr(lr*1e6,2)-47.009*lr*1e6+4.7061)*wr*1e6+(-74.026*pwr(lr*1e6,2)+47.818*lr*1e6-4.9076)))*1e-15, 1e-18)'
+Rsub1_rf     = 'max(((-173.25*lr*1e6+30.089)*pwr(wr*1e6,2)+(1110*lr*1e6-81.61)*wr*1e6+(-7105.6*lr*1e6+1996.8))*pwr(nf,1.7573*lr*1e6-0.8936), 1e-3)'
+Rsub2_rf     = 'max(((-2.52*lr*1e6+0.4097)*pwr(wr*1e6,2)+(16.422*lr*1e6-2.5923)*wr*1e6+(-21.611*lr*1e6+2.9913))*nf+((43.175*lr*1e6-5.3693)*pwr(wr*1e6,2)+(-232.18*lr*1e6+24.958)*wr*1e6+(399*lr*1e6+31.75)), 1e-3)'
+Rsub3_rf     = 'max(((-318.02*lr*1e6+94.625)*pwr(wr*1e6,2)+(4878.4*lr*1e6-1449.3)*wr*1e6+(-18771*lr*1e6+5701.4))+((1288.3*lr*1e6-389.18)*pwr(wr*1e6,2)+(-18714*lr*1e6+5649.5)*wr*1e6+(59353*lr*1e6-18005))/NF, 1e-3)'
+Djdb_AREA_rf = 'nf/2*wr*(0.8-0.14)*1e-6'
+Djdb_PJ_rf   = '(1+1.2547e-7/wr)*nf*wr'
+Djsb_AREA_rf = 'wr*(0.8-0.07)*2*1e-6+(nf/2-1)*wr*(0.8-0.14)*1e-6'
+Djsb_PJ_rf   = '(1+1.2547e-7/wr)*nf*wr'
+Rdc_n18      = 'max((0.1008/(wr*1e6)+0.102*nf), 1e-3)'
+Rsc_n18      = 'max((0.1008/(wr*1e6)+0.102*nf), 1e-3)'   
+Cgdo_n18     = 'max((0+dcgdo_n18_rf), 0)'
+Cgso_n18     = 'max((0+dcgso_n18_rf), 0)'
+Cj_n18       = 'max((0+dcj_n18_rf), 0)'
+Cjsw_n18     = 'max((0+dcjsw_n18_rf), 0)'
+Pvag_n18     = '-((0.0733*lr*1000000-0.0117)*pwr(wr*1000000,2)+(-1.02*lr*1000000+0.1431)*wr*1000000+(3.3992*lr*1000000-0.2917))*pwr(nf,(0.0508*lr*1000000-0.0097)*pwr(wr*1000000,2)+(-0.3633*lr*1000000+0.1088)*wr*1000000+(-0.24*lr*1000000+0.0165))'
*****************************************
Lgate       2 20  1p
Rgate       20 21 Rg_rf
Cgd_ext     20 11 Cgd_rf
Cgs_ext     20 31 Cgs_rf
Cds_ext     15 31 Cds_rf
Rds         11 15 0.01
Ldrain       1 11 1p
Lsource      3 31 1p
*****************************************
Djdb  12 11
+ ndio18_rf
+ AREA  = Djdb_AREA_rf
+ PJ    = Djdb_PJ_rf 
***
Djsb  32 31
+ ndio18_rf
+ AREA  = Djsb_AREA_rf
+ PJ    = Djsb_PJ_rf
*****************************************
Rsub1      41  4  Rsub1_rf
Rsub2      41  12 Rsub2_rf
Rsub3      41  32 Rsub3_rf
*
* --------- ideal mos transistor ----------------------
MAIN 11 21 31 41 n18_rf L=lr W=wr m=nf AD = 0 AS = 0 PD = 0 PS = 0
* MOS Model
.model  n18_rf  nmos
+level = 49
**************************************************************
*               MODEL FLAG PARAMETERS 
**************************************************************
+lmin    = 1.6e-007        lmax    = 1.2e-006        wmin    = 4.8e-007      
+wmax    = 1.002e-005      version = 3.24             mobmod  = 1             
+capmod  = 3               nqsmod  = 0               binunit = 2             
**************************************************************
*               GENERAL MODEL PARAMETERS 
**************************************************************
+tref    = 25              xl      = '1.8e-008+DXL_N18_RF'        xw      = '0+DXW_N18_RF'             
+tox     = '3.87e-009+DTOX_N18_RF'        toxm    = 3.87e-009       wint    = -1.4450482E-09      
+lint    = 1.5757085E-08     dlc     = 8.5e-009        dwc     = 4.5e-008      
+hdif    = 2e-007          ldif    = 7e-008          ll      = 2.6352781e-016
+wl      = -2.3664573e-016  lln     = 1.1205959       wln     = 1.0599999     
+lw      = -2.2625584e-016  ww      = -3.640969e-014  lwn     = 0.92          
+wwn     = 0.8768474       lwl     = -2.0576711e-022  wwl     = -4e-021       
+cgso    = 'Cgso_n18'               cgdo    = 'Cgdo_n18'               xpart   = 1   
+rdc ='Rdc_n18' rsc='Rsc_n18'          
**************************************************************
*               EXPERT PARAMETERS 
**************************************************************
+vth0    = '0.39+DVTH_N18_RF'        wvth0   = -2.9709472e-008  pvth0   = '5e-016+DPVTH0_N18_RF'                
+k1      = 0.6801043       wk1     = -2.489684e-008  pk1     = 1.3e-015      
+k2      = -0.049978       k3      = 10              k3b     = -3            
+nlx     = 7.545103e-008   dvt0    = 1.3             dvt1    = 0.5771635     
+dvt2    = -0.1717554      dvt0w   = 0               dvt1w   = 0             
+dvt2w   = 0               nch     = 3.8694e+017     voff    = -0.103        
+lvoff   = -3.3e-009       nfactor = 1.25            lnfactor= 4.5e-008      
+cdsc    = 0               cdscb   = 0               cdscd   = 0.0001        
+cit     = 0               u0      = 0.032953        lu0     = 2.3057663e-011
+wu0     = -3.1009695e-009  ua      = -1.03e-009      lua     = 7.734979e-019 
+pua     = -1e-024         ub      = 2.3667e-018     uc      = 1.2e-010      
+puc     = 1.5e-024        xj      = 1.6e-007        w0      = 5.582015e-007 
+prwg    = 0.4             prwb    = -0.24           wr      = 1             
+rdsw    = 55.54972        a0      = 0.83            ags     = 0.32          
+a1      = 0               a2      = 0.99            b0      = 6e-008        
+b1      = 0               vsat    = 82500           pvsat   = -8.3e-010     
+keta    = -0.003          lketa   = -1.7e-009       dwg     = -5.96e-009    
+dwb     = 4.5e-009        alpha0  = 1.7753978e-008  beta0   = 11.168394     
+pclm    = 1.2             ppclm   = 2.9999999e-015  pdiblc1 = 0.025         
+pdiblc2 = 0.0038          ppdiblc2= 2.7000001e-016  pdiblcb = 0             
+drout   = 0.56            pvag    = 'Pvag_n18'               pscbe1  = 3.45e+008     
+pscbe2  = 1e-006          delta   = 0.01            eta0    = 0.028000001   
+etab    = -0.027000001    dsub    = 0.4             elm     = 5             
+alpha1  = 0.1764          lalpha1 = 7.625e-009    
**************************************************************
*               CAPACITANCE PARAMETERS 
**************************************************************
+cf      = 0               acde    = 0.64            moin    = 24            
+noff    = 1.2025        CJ       = 'Cj_n18'
+CJSW     = 'Cjsw_n18'   CGBO=0

**************************************************************
*               TEMPERATURE PARAMETERS 
**************************************************************
+kt1     = -0.2572866      kt1l    = -1e-009         kt2     = -0.04         
+ute     = -1.55           ua1     = 1.76e-009       lua1    = 6e-018        
+wua1    = -1.1e-016       pua1    = -5e-025         ub1     = -2.4e-018     
+uc1     = -1e-010         luc1    = 1.6999999e-017  puc1    = -3e-024       
+prt     = -55             at      = 37000           pat     = -7.5e-010     
**************************************************************
*               NOISE PARAMETERS 
**************************************************************
+NOIMOD   = 2                   NOIA     = 8.2282E+19            NOIB     = 1.3327E+04    
+NOIC     = -2.4937E-14         EM       = 1.7767E+07            EF       = 8.1800E-01 
**************************************************************
.model ndio18_rf D
+LEVEL    = 3                   JS       = 3.52e-07            JSW      = 1e-15            
+N        = 1.0233              IK       = 1.52e+05            
+IKR      = 2.78e+05            BV       = 11.0                IBV      = 277.78              
+TRS      = 1.51e-03            EG       = 1.16                TREF     = 25.0                
+XTI      = 3.0                             
+CJ       = 9.68E-04
+CJSW     = 4.18E-10
+RS       = 8.89e-09
+MJ       = 0.346               PB       = 0.7                 MJSW     = 0.538               
+PHP      = 1                   CTA      = 0.000842            CTP      = 0.000669            
+TPB      = 0.00147             TPHP     = 0.000868            TLEV     = 1
+TLEVC    = 1                   FC       = 0                   FCS      = 0 
.ends n18_ckt_rf
***************************
* 1.8V RF DNWMOS Subcircuit
***************************
* 11=drain, 2=gate, 31=source, 4=bulk, 5=DNW
* lr=gate length, wr=finger width, nf=finger number, laddr=DNW diode add length, waddr=DNW diode add width
.subckt dnw18_ckt_rf 1 2 3 4 5 lr=l wr=w nf=finger laddr=ladd waddr=wadd
* scalable unit parameter
* euqivalent circuit saclable parameter
.param
+Rg_rf        = 'max(((724.84*pwr(lr*1e6,2)-356.18*lr*1e6+50.477)+(-72.591*pwr(lr*1e6,2)+34.823*lr*1e6-4.3737)*wr*1e6+(-709.9*pwr(lr*1e6,2)+340.42*lr*1e6-49.734)/(wr*1e6))+((-5161.5*pwr(lr*1e6,2)+1999.2*lr*1e6-33.119)+(531.35*pwr(lr*1e6,2)-224.13*lr*1e6+12.828)*wr*1e6+(3902.6*pwr(lr*1e6,2)-164.08*lr*1e6+386.39)/(wr*1e6))/nf,1e-3)'
+Cgd_rf       = 'max((((0.6677*pwr(lr*1e6,2)-0.4222*lr*1e6+0.0529)*pwr(wr*1e6,2)+(-5.7464*pwr(lr*1e6,2)+3.8016*lr*1e6-0.1298)*wr*1e6+(3.275*pwr(lr*1e6,2)-2.272*lr*1e6+0.6075))*nf+((-3.5823*pwr(lr*1e6,2)+2.4353*lr*1e6-0.3546)*pwr(wr*1e6,2)+(30.068*pwr(lr*1e6,2)-20.101*lr*1e6+2.8423)*wr*1e6+(-23.613*pwr(lr*1e6,2)+15.794*lr*1e6-1.9974)))*1e-15, 1e-18)'
+Cgs_rf       = 'max((((0.0651*pwr(lr*1e6,2)-0.0346*lr*1e6+0.004)*pwr(wr*1e6,2)+(-0.701*pwr(lr*1e6,2)+0.3523*lr*1e6-0.0371)*wr*1e6+(1.0807*pwr(lr*1e6,2)-0.5396*lr*1e6+0.061))*pwr(nf,2)+((-0.1448*pwr(lr*1e6,2)-0.1172*lr*1e6+0.0525)*pwr(wr*1e6,2)+(1.1016*pwr(lr*1e6,2)+2.1538*lr*1e6-0.8227)*wr*1e6+(-11.232*pwr(lr*1e6,2)+1.8929*lr*1e6+0.7917))*nf+((-2.1156*pwr(lr*1e6,2)+2.368*lr*1e6-0.5178)*pwr(wr*1e6,2)+(33.552*pwr(lr*1e6,2)-34.449*lr*1e6+6.9433)*wr*1e6+(-54.224*pwr(lr*1e6,2)+52.226*lr*1e6-7.2535)))*1e-15, 1e-18)'
*+Cgs_rf       = 'max((((-2.4185E-18*lr*1e6*lr*1e6+1.9748E-18*lr*1e6-1.1477E-19)*wr*1e6*wr*1e6+(1.7561E-17*lr*1e6*lr*1e6-1.5834E-17*lr*1e6+3.0446E-18)*wr*1e6+(5.1244E-17*lr*1e6*lr*1e6-1.8280E-17*lr*1e6+2.1420E-18))*nf*nf+((2.3832E-16*lr*1e6*lr*1e6-1.9105E-16*lr*1e6+3.0968E-17)*wr*1e6*wr*1e6+(-1.5807E-15*lr*1e6*lr*1e6+1.3096E-15*lr*1e6-2.9961E-16)*wr*1e6+(-3.3719E-15*lr*1e6*lr*1e6+2.8975E-15*lr*1e6+3.0622E-16))*nf+((2.8363e-16*lr*1e6*lr*1e6-1.128E-16*lr*1e6+3.4224E-17)*wr*1e6*wr*1e6+(-6.1212e-15*lr*1e6*lr*1e6+2.5933E-15*lr*1e6-7.0304e-16)*wr*1e6+(3.4536E-14*lr*1e6*lr*1e6-1.4597E-14*lr*1e6+4.3951E-15))), 1e-18)'
+Cds_rf       = 'max((((1.2656*pwr(lr*1e6,2)-0.8625*lr*1e6+0.1269)*pwr(wr*1e6,2)+(-14.055*pwr(lr*1e6,2)+8.8032*lr*1e6-0.7362)*wr*1e6+(16.189*pwr(lr*1e6,2)-11.156*lr*1e6+1.6503))*nf+((-6.6026*pwr(lr*1e6,2)+3.9526*lr*1e6-0.3798)*pwr(wr*1e6,2)+(76.57*pwr(lr*1e6,2)-47.009*lr*1e6+4.7061)*wr*1e6+(-74.026*pwr(lr*1e6,2)+47.818*lr*1e6-4.9076)))*1e-15, 1e-18)'
+Rsub1_rf     = 'max(((-173.25*lr*1e6+30.089)*pwr(wr*1e6,2)+(1110*lr*1e6-81.61)*wr*1e6+(-7105.6*lr*1e6+1996.8))*pwr(nf,1.7573*lr*1e6-0.8936), 1e-3)'
+Rsub2_rf     = 'max(((-2.52*lr*1e6+0.4097)*pwr(wr*1e6,2)+(16.422*lr*1e6-2.5923)*wr*1e6+(-21.611*lr*1e6+2.9913))*nf+((43.175*lr*1e6-5.3693)*pwr(wr*1e6,2)+(-232.18*lr*1e6+24.958)*wr*1e6+(399*lr*1e6+31.75)), 1e-3)'
+Rsub3_rf     = 'max(((-318.02*lr*1e6+94.625)*pwr(wr*1e6,2)+(4878.4*lr*1e6-1449.3)*wr*1e6+(-18771*lr*1e6+5701.4))+((1288.3*lr*1e6-389.18)*pwr(wr*1e6,2)+(-18714*lr*1e6+5649.5)*wr*1e6+(59353*lr*1e6-18005))/NF, 1e-3)'
+Djdb_AREA_rf = 'nf/2*wr*(0.8-0.14)*1e-6'
+Djdb_PJ_rf   = '(1+1.2547e-7/wr)*nf*wr'
+Djsb_AREA_rf = 'wr*(0.8-0.07)*2*1e-6+(nf/2-1)*wr*(0.8-0.14)*1e-6'
+Djsb_PJ_rf   = '(1+1.2547e-7/wr)*nf*wr'
+Djbdn_AREA_rf= '(2*0.8*1e-6+lr*nf+0.8*1e-6*(nf-1)+2*laddr)*(wr+2*waddr)'
+Djbdn_PJ_rf  = '2*(2*0.8*1e-6+lr*nf+0.8*1e-6*(nf-1)+wr+2*(laddr+waddr))'
+Rdc_n18      = 'max((0.1008/(wr*1e6)+0.102*nf), 1e-3)' 
+Rsc_n18      = 'max((0.1008/(wr*1e6)+0.102*nf), 1e-3)' 
+Cgdo_n18     = 'max((0+dcgdo_n18_rf), 0)'
+Cgso_n18     = 'max((0+dcgso_n18_rf), 0)'
*+Cf_n18       = 'max((0+dcf_n18_rf), 0)'
*+Cgdl_n18     = 'max((0+dcgdl_n18_rf), 0)'
*+Cgsl_n18     = 'max((0+dcgsl_n18_rf), 0)'
+Cj_n18       = 'max((0+dcj_n18_rf), 0)'
+Cjsw_n18     = 'max((0+dcjsw_n18_rf), 0)'
*+Cjswg_n18    = 'max((0+dcjswg_n18_rf), 0)'
+Pvag_n18     = '-((0.0733*lr*1000000-0.0117)*pwr(wr*1000000,2)+(-1.02*lr*1000000+0.1431)*wr*1000000+(3.3992*lr*1000000-0.2917))*pwr(nf,(0.0508*lr*1000000-0.0097)*pwr(wr*1000000,2)+(-0.3633*lr*1000000+0.1088)*wr*1000000+(-0.24*lr*1000000+0.0165))'
*****************************************
Lgate       2 20  1p
Rgate       20 21 Rg_rf
Cgd_ext     20 11 Cgd_rf
Cgs_ext     20 31 Cgs_rf
Cds_ext     15 31 Cds_rf
Rds         11 15 0.01
Ldrain       1 11 1p
Lsource      3 31 1p
*****************************************
Djdb  12 11
+ ndio18_rf
+ AREA  = Djdb_AREA_rf
+ PJ    = Djdb_PJ_rf 
***
Djsb  32 31
+ ndio18_rf
+ AREA  = Djsb_AREA_rf
+ PJ    = Djsb_PJ_rf
***
Djbdn  4 5
+ diobpw_rf
+ AREA  = Djbdn_AREA_rf
+ PJ    = Djbdn_PJ_rf
*****************************************
Rsub1      41  4  Rsub1_rf
Rsub2      41  12 Rsub2_rf
Rsub3      41  32 Rsub3_rf
*
* --------- ideal mos transistor ----------------------
MAIN 11 21 31 41 dnw18_rf L=lr W=wr m=nf AD = 0 AS = 0 PD = 0 PS = 0
* MOS Model
.MODEL dnw18_rf NMOS
+LEVEL = 49
**************************************************************
*               MODEL FLAG PARAMETERS 
**************************************************************
+lmin    = 1.6e-007        lmax    = 1.2e-006        wmin    = 4.8e-007      
+wmax    = 1.002e-005      version = 3.24             mobmod  = 1             
+capmod  = 3               nqsmod  = 0               binunit = 2             
**************************************************************
*               GENERAL MODEL PARAMETERS 
**************************************************************
+tref    = 25              xl      = '1.8e-008+DXL_N18_RF'        xw      = '0+DXW_N18_RF'             
+tox     = '3.87e-009+DTOX_N18_RF'        toxm    = 3.87e-009       wint    = -1.4450482E-09      
+lint    = 1.5757085E-08     dlc     = 8.5e-009        dwc     = 4.5e-008      
+hdif    = 2e-007          ldif    = 7e-008          ll      = 2.6352781e-016
+wl      = -2.3664573e-016  lln     = 1.1205959       wln     = 1.0599999     
+lw      = -2.2625584e-016  ww      = -3.640969e-014  lwn     = 0.92          
+wwn     = 0.8768474       lwl     = -2.0576711e-022  wwl     = -4e-021       
+cgso    = 'Cgso_n18'               cgdo    = 'Cgdo_n18'               xpart   = 1   
+rdc ='Rdc_n18' rsc='Rsc_n18'          
**************************************************************
*               EXPERT PARAMETERS 
**************************************************************
+vth0    = '0.39+DVTH_N18_RF'        wvth0   = -2.9709472e-008  pvth0   = '5e-016+DPVTH0_N18_RF'                
+k1      = 0.6801043       wk1     = -2.489684e-008  pk1     = 1.3e-015      
+k2      = -0.049978       k3      = 10              k3b     = -3            
+nlx     = 7.545103e-008   dvt0    = 1.3             dvt1    = 0.5771635     
+dvt2    = -0.1717554      dvt0w   = 0               dvt1w   = 0             
+dvt2w   = 0               nch     = 3.8694e+017     voff    = -0.103        
+lvoff   = -3.3e-009       nfactor = 1.25            lnfactor= 4.5e-008      
+cdsc    = 0               cdscb   = 0               cdscd   = 0.0001        
+cit     = 0               u0      = 0.032953        lu0     = 2.3057663e-011
+wu0     = -3.1009695e-009  ua      = -1.03e-009      lua     = 7.734979e-019 
+pua     = -1e-024         ub      = 2.3667e-018     uc      = 1.2e-010      
+puc     = 1.5e-024        xj      = 1.6e-007        w0      = 5.582015e-007 
+prwg    = 0.4             prwb    = -0.24           wr      = 1             
+rdsw    = 55.54972        a0      = 0.83            ags     = 0.32          
+a1      = 0               a2      = 0.99            b0      = 6e-008        
+b1      = 0               vsat    = 82500           pvsat   = -8.3e-010     
+keta    = -0.003          lketa   = -1.7e-009       dwg     = -5.96e-009    
+dwb     = 4.5e-009        alpha0  = 1.7753978e-008  beta0   = 11.168394     
+pclm    = 1.2             ppclm   = 2.9999999e-015  pdiblc1 = 0.025         
+pdiblc2 = 0.0038          ppdiblc2= 2.7000001e-016  pdiblcb = 0             
+drout   = 0.56            pvag    = 'Pvag_n18'               pscbe1  = 3.45e+008     
+pscbe2  = 1e-006          delta   = 0.01            eta0    = 0.028000001   
+etab    = -0.027000001    dsub    = 0.4             elm     = 5             
+alpha1  = 0.1764          lalpha1 = 7.625e-009    
**************************************************************
*               CAPACITANCE PARAMETERS 
**************************************************************
+cf      = 0               acde    = 0.64            moin    = 24            
+noff    = 1.2025        CJ       = 'Cj_n18'
+CJSW     = 'Cjsw_n18'           CGBO=0

**************************************************************
*               TEMPERATURE PARAMETERS 
**************************************************************
+kt1     = -0.2572866      kt1l    = -1e-009         kt2     = -0.04         
+ute     = -1.55           ua1     = 1.76e-009       lua1    = 6e-018        
+wua1    = -1.1e-016       pua1    = -5e-025         ub1     = -2.4e-018     
+uc1     = -1e-010         luc1    = 1.6999999e-017  puc1    = -3e-024       
+prt     = -55             at      = 37000           pat     = -7.5e-010     
**************************************************************
*               NOISE PARAMETERS 
**************************************************************
+NOIMOD   = 2                   NOIA     = 8.2282E+19            NOIB     = 1.3327E+04    
+NOIC     = -2.4937E-14         EM       = 1.7767E+07            EF       = 8.1800E-01 
**************************************************************
.model ndio18_rf D
+LEVEL    = 3                   JS       = 3.52e-07            JSW      = 1e-15            
+N        = 1.0233              IK       = 1.52e+05            
+IKR      = 2.78e+05            BV       = 11.0                IBV      = 277.78              
+TRS      = 1.51e-03            EG       = 1.16                TREF     = 25.0                
+XTI      = 3.0                             
+CJ       = 9.68E-04
+CJSW     = 4.18E-10
+RS       = 8.89e-09
+MJ       = 0.346               PB       = 0.7                 MJSW     = 0.538               
+PHP      = 1                   CTA      = 0.000842            CTP      = 0.000669            
+TPB      = 0.00147             TPHP     = 0.000868            TLEV     = 1
+TLEVC    = 1                   FC       = 0                   FCS      = 0 
.model diobpw_rf D 
*   
+LEVEL    = 3                   JS       = 1.50E-07            JSW      = 1.00E-15            
+N        = 1.0213              RS       = 2.51E-08            IK       = 2.40E+05            
+IKR      = 1.04E+05            BV       = 15.0                IBV      = 1.04E+02                
+TRS      = 1.77E-03            CTA      = 0.0012              CTP      = 0.00107                
+EG       = 1.16                TREF     = 25.0                TPB      = 0.0019               
+TPHP     = 0.00193             XTI      = 3.0                 CJ       = 0.000536            
+MJ       = 0.343               PB       = 0.693               CJSW     = 3.22E-10            
+MJSW     = 0.361               PHP      = 0.715               TLEV     = 1
+TLEVC    = 1      		AREA     = 9.6E-9              PJ       = 4E-4  
+FC       = 0                   FCS      = 0
.ends dnw18_ckt_rf
*************************
* 1.8V RF PMOS Subcircuit
*************************
* 11=drain, 2=gate, 31=source, 4=bulk
* lr=gate length, wr=finger width, nf=finger number
.subckt p18_ckt_rf 1 2 3 4 lr=l wr=w nf=finger
* scalable unit parameter
* euqivalent circuit saclable parameter
.param
+Cgs_rf    = 'max((((6.2506e-17*lr*lr*1e6*1e6-2.9036e-17*lr*1e6+3.9433e-18)*exp((-2.0989*lr*lr*1e6*1e6+8.7703e-1*lr*1e6+2.6579e-1)*wr*1e6))*nf*nf+((4.4788e-16*lr*lr*1e6*1e6-4.0771e-16*lr*1e6-1.0686e-17)*wr*1e6+(-2.3431e-15*lr*lr*1e6*1e6+2.2217e-15*lr*1e6+3.6221e-16))*nf+((6.7052e-15*lr*lr*1e6*1e6-6.2642e-15*lr*1e6+2.7578e-16)*log(wr*1e6)+(-1.2255e-14*lr*lr*1e6*1e6+1.562e-14*lr*1e6-1.487e-16))), 1e-18)'
+Rg_rf        = 'max((((17236*lr*lr*1e6*1e6+181.46*lr*1e6+149.85)*pwr(wr*1e6,(1.3797*lr*lr*1e6*1e6-2.4198*lr*1e6-0.48)))*pwr(nf,(0.5573*lr*lr*1e6*1e6-0.1633*lr*1e6+0.1623)*log(wr*1e6)+(-1.0151*lr*lr*1e6*1e6-0.1544*lr*1e6-0.981))), 1e-3)'
+Rsub1_rf     = 'max((0.0023528*nf*nf-0.56425*nf+61.816), 1e-3)'
+Rsub2_rf     = 'max((-11.603*log(nf)+72.058), 1e-3)'
+Rsub3_rf     = 'max((-1065.3*log(nf)+5768.9), 1e-3)'
+Cgd_rf       = 'max((((5.375E-17*lr*lr*1e6*1e6-1.08E-17*lr*1e6+4.4E-16)*wr*1e6+(-3.9974E-16*lr*lr*1e6*1e6+6.9454E-16*lr*1e6+(1.3021E-16*lr*lr*1e6*1e6+2.0833E-17*lr*1e6+9.2031E-17)))*nf+(1.7802E-17*wr*wr*1e6*1e6-3.4928E-16*wr*1e6+6.1859E-16)), 1e-18)'
+Cds_rf       = 'max(((4.1455e-16*lr*lr*1e6*1e6-3.5118e-16*lr*1e6+6.4154e-17)*wr*wr*1e6*1e6+(-9.4276e-16*lr*lr*1e6*1e6+8.0336e-16*lr*1e6+1.1269e-16)*wr*1e6+(-4.1859e-16*lr*lr*1e6*1e6+9.8925e-17*lr*1e6+2.1732e-16))*nf+((-4.9953e-17*lr*1e6*lr*1e6+1.011e-16*lr*1e6+5.9634e-17)*wr*1e6+(-1.7041e-15*lr*lr*1e6*1e6+1.571e-15*lr*1e6+4.9801e-16)), 1e-18)'
+Djdb_AREA_rf = '(nf/2*(0.8-2*0.07)*wr)*1e-6'
+Djdb_PJ_rf   = '(1+1.287e-7/wr)*nf*wr'
+Djsb_AREA_rf = '((nf/2-1)*(0.8-2*0.07)*wr+(0.8-0.07)*wr*2)*1e-6'
+Djsb_PJ_rf   = '(1+1.287e-7/wr)*nf*wr'
+Cgdo_p18_rf     = 'max((0+dcgdo_p18_rf), 0)'
+Cgso_p18_rf     = 'max((0+dcgso_p18_rf), 0)'
+Cj_p18_rf    = 'max((0+dcj_p18_rf), 0)'
+Cjsw_p18_rf     = 'max((0+dcjsw_p18_rf), 0)'
+Rdc_p18_rf       = 'max((32.428*exp(-0.3464*wr*1e6))*pwr(nf, 0.1502*exp(0.1353*wr*1e6)), 1e-3)'
+Rsc_p18_rf       = 'max((32.428*exp(-0.3464*wr*1e6))*pwr(nf, 0.1502*exp(0.1353*wr*1e6)), 1e-3)'
*****************************************
Lgate       2 20  1p
Rgate       20 21 Rg_rf
Cgd_ext     20 11 Cgd_rf
Cgs_ext     20 31 Cgs_rf
Cds_ext     15 31 Cds_rf
Rds         11 15 0.01
Ldrain       1 11 1p
Lsource      3 31 1p
*****************************************
Djdb  11 12
+ pdio18_rf
+ AREA  = Djdb_AREA_rf
+ PJ    = Djdb_PJ_rf 
***
Djsb  31 32
+ pdio18_rf
+ AREA  = Djsb_AREA_rf
+ PJ    = Djsb_PJ_rf
*****************************************
Rsub1      41  4  Rsub1_rf
Rsub2      41  12 Rsub2_rf
Rsub3      41  32 Rsub3_rf
*
* --------- ideal mos transistor ----------------------
MAIN 11 21 31 41 p18_rf L=lr W=wr m=nf AD = 0 AS = 0 PD = 0 PS = 0
* MOS Model
.MODEL p18_rf PMOS
+LEVEL = 49
*
* GENERAL PARAMETERS
*
+CALCACM  = 1
+LMIN     = 1.6E-7              LMAX     = 5.2E-7              WMIN     = 4.8E-7              
+WMAX     = 1.002E-5            TNOM     = 25.0                VERSION  = 3.24                 
+TOX      = '3.74E-09+DTOX_P18_RF'  TOXM     = 3.74E-09            XJ       = 1.7000001E-07       
+NCH      = 5.5000000E+17       LLN      = 1.0000000           LWN      = 1.0000000           
+WLN      = 1.0450000           WWN      = 1.0000000           LINT     = 1.3800000E-08       
+LL       = 3.4000000E-15       LW       = -3.3600000E-16      LWL      = 0.00                
+WINT     = -5.0000000E-09       WL       = 3.5904200E-15       WW       = -1.8999999E-15      
+WWL      = -1.1205000E-21      MOBMOD   = 1                   BINUNIT  = 2                   
+XL       = '-5.7E-09+DXL_P18_RF'   XW       = '0.00+DXW_P18_RF'      DWG      = -1.7361970E-08          
+DWB      = 2.0000000E-08       
* DIODE PARAMETERS
+ACM      = 12                  LDIF     = 7.00E-08            HDIF     = 2.00E-07            
+RSH      = 7.83                RD       = 0                   RS       = 0                   
+RSC      = 'Rsc_p18_rf'               RDC      = 'Rdc_p18_rf'                 
*
* THRESHOLD VOLTAGE PARAMETERS
*
+VTH0     = '-0.41+DVTH_P18_RF'   WVTH0    = 1.2675420E-08       PVTH0    = '-1.2500000E-15+DPVTH0_P18_RF'     
+K1       = 0.5872390           LK1      = 3.5532110E-09       K2       = 7.0906860E-03       
+K3       = 2.5999999           DVT0     = 0.7194931           DVT1     = 0.2467441           
+DVT2     = 7.8089680E-02       DVT0W    = 0.00                DVT1W    = 8.0000000E+05       
+DVT2W    = 0.00                NLX      = 9.0000000E-08       W0       = 0.00                
+K3B      = 2.4862001           NGATE    = 3.1680000E+20               
*
* MOBILITY PARAMETERS
*
+VSAT     = 1.0000000E+05       UA       = 2.8500000E-10       LUA      = 5.5000000E-18       
+PUA      = -2.0000000E-24      UB       = 1.0000000E-18       UC       = -4.7700000E-11      
+WUC      = 3.1668000E-17       PUC      = -2.5000000E-24      RDSW     = 4.5500000E+02       
+PRWB     = -0.4000000          PRWG     = 0.00                WR       = 1.0000000           
+U0       = 8.6610000E-03       LU0      = -2.0000000E-11      WU0      = 1.3815350E-10       
+A0       = 1.0000000           KETA     = 2.0000000E-02       LKETA    = -8.5000000E-09      
+PKETA    = 5.0000000E-16       A1       = 0.00                A2       = 0.9900000           
+AGS      = 0.2000000           B0       = 6.3000000E-08       B1       = 0.00                
*
* SUBTHRESHOLD CURRENT PARAMETERS
*
+VOFF     = -9.5000000E-02      LVOFF    = -1.7000000E-09      WVOFF    = -1.9999999E-09      
+PVOFF    = -1.0000000E-16      NFACTOR  = 0.9000000           LNFACTOR = 1.0000000E-07       
+PNFACTOR = -5.0000000E-15      CIT      = 0.00                CDSC     = 0.00                
+CDSCB    = 0.00                CDSCD    = 0.00                ETA0     = 4.0000000E-02       
+ETAB     = -2.5000000E-02      DSUB     = 0.5600000           
*
* ROUT PARAMETERS
*
+PCLM     = 0.7000000           PDIBLC1  = 0.00                PDIBLC2  = 7.0000000E-03       
+PDIBLCB  = 0.00                DROUT    = 0.5600000           PSCBE1   = 4.0000000E+08       
+PSCBE2   = 1.0000000E-07       PVAG     = 0.00                DELTA    = 1.0000000E-02       
+ALPHA0   = 7.0000000E-08       ALPHA1   = 7.0491700           BETA0    = 22.8424000          
+LBETA0   = -7.5000000E-08         
*
* TEMPERATURE EFFECTS PARAMETERS
*
+KT1      = -0.2577007          KT2      = -3.0979900E-02      LKT2     = -3.0000000E-09      
+PKT2     = -6.5331750E-16      AT       = 1.0000000E+04       PAT      = -1.0000000E-09      
+UTE      = -1.2703574          UA1      = 5.3866300E-10       WUA1     = 1.1000000E-16       
+PUA1     = -2.3700001E-24      UB1      = -2.0709999E-18      UC1      = 2.0609721E-11       
+KT1L     = -8.0000000E-09      PRT      = 90.0000000          
*
* CAPACITANCE PARAMETERS
*
+CJ       = 'Cj_p18_rf'                   MJ       = 0.415               PB       = 0.817                   
+CJSW     = 'Cjsw_p18_rf'                    MJSW     = 0.489               PBSW     = 1               
+CJSWG    = 0                   MJSWG    = 0.489               PBSWG    = 1       
+TPB      = 0.00153             TPBSW    = 0.00117             TPBSWG   = 0.00117
+TCJ      = 0.000876            TCJSW    = 0.000745            TCJSWG   = 0.000745
+JS       = 1.66E-07            JSW      = 1.2E-13             NJ       = 1.0384   
+XTI      = 4.5                 NQSMOD   = 0                   ELM      = 5 
+CGDO     = 'Cgdo_p18_rf'        CGSO     = 'Cgso_p18_rf'   CGBO = 0       TLEVC    = 1            
+CAPMOD   = 3                   XPART    = 1                   CF       = 0.00                                    
+ACDE     = 0.8505076           MOIN     = 14.95341            NOFF     = 1.431824              
+DLC      = -1.5E-09
*
* NOISE PARAMETERS
*
+NOIMOD   = 2                   NOIA     = 3.3617E+18            NOIB     = 1.9536E+05    
+NOIC     = 5.2658E-12          EM       = 6.2548E+07            EF       = 1.1307E+00 
*
* Diode Model 
.model pdio18_rf d
*
+LEVEL    = 3                   JS       = 1.66E-07            JSW      = 1E-15             
+N        = 1.0135              RS       = 8.77E-09            IK       = 4.03E+05            
+IKR      = 2.78E+05            BV       = 11.0                IBV      = 277.78              
+TRS      = 1.78E-03            EG       = 1.16                TREF     = 25.0                
+XTI      = 3.0                 CJ       = 0.00107             MJ       = 0.415               
+PB       = 0.817               CJSW     = 5.07E-10            MJSW     = 0.489               
+PHP      = 0.95                CTA      = 0.000876            CTP      = 0.000745            
+TPB      = 0.00153             TPHP      = 0.00117            TLEV     = 1
+TLEVC    = 1            FC       = 0                   FCS      = 0   
.ends p18_ckt_rf
*************************
* 3.3V RF NMOS Subcircuit
*************************
* 11=drain, 2=gate, 31=source, 4=bulk
* lr=gate length, wr=finger width, nf=finger number
.subckt n33_ckt_rf 1 2 3 4 lr=l wr=w nf=finger
* scalable unit parameter
* euqivalent circuit saclable parameter
.param
+Rg_rf        = 'max((((337.44*lr*lr*1e6*1e6-636.15*lr*1e6+1247.8)*pwr(wr*1e6,(0.0345*lr*lr*1e6*1e6-0.0673*lr*1e6-0.8144)))*pwr(nf,(0.01549*lr*lr*1e6*1e6-0.02983*lr*1e6+0.10754)*log(wr*1e6)+(-0.01723*lr*lr*1e6*1e6+0.03465*lr*1e6-0.95262))),1e-3)'
+Cgd_rf       = 'max((((-1.019487e-18*lr*lr*1e6*1e6+2.093231E-18*lr*1e6-5.621744E-18)*wr*wr*1e6*1e6+(-7.0297E-17*lr*lr*1e6*1e6+1.4369E-16*lr*1e6+3.8644E-16)*wr*1e6+(9.4974E-18*lr*lr*1e6*1e6+3.9394E-17*lr*1e6+2.3454E-16))*nf+((-4.8156E-18*lr*lr*1e6*1e6+1.1596E-16*lr*1e6-2.1673E-17)*wr*wr*1e6*1e6+(4.816E-16*lr*lr*1e6*1e6-1.2046E-15*lr*1e6+8.1E-19)*wr*1e6+(-1.5056E-16*lr*lr*1e6*1e6+7.2245E-16*lr*1e6+2.1267E-16))),1e-18)'
+Cgs_rf       = 'max(((-1.7423e-17*lr*lr*1e6*1e6+3.3616E-17*lr*1e6+7.4972E-19)*wr*wr*1e6*1e6+(-8.3169E-17*lr*lr*1e6*1e6+2.8529E-16*lr*1e6+2.5325E-16)*wr*1e6+(-5.1487E-16*lr*lr*1e6*1e6+9.9831E-16*lr*1e6+3.2256E-16))*nf+((-2.5956E-17*lr*lr*1e6*1e6-2.5684E-17*lr*1e6+1.5362E-16)*wr*wr*1e6*1e6+(-3.6262E-15*lr*lr*1e6*1e6+6.3722E-15*lr*1e6-3.7861E-15)*wr*1e6+(8.4615E-15*lr*lr*1e6*1e6-1.4192E-14*lr*1e6+7.9308E-15)),1e-18)'
+Cds_rf       = 'max(((-8.3173e-17*lr*lr*1e6*1e6+1.4664E-16*lr*1e6-3.1474E-17)*wr*wr*1e6*1e6+(4.9488E-16*lr*lr*1e6*1e6-8.6038E-16*lr*1e6+4.8447E-16)*wr*1e6+(-6.5021E-16*lr*lr*1e6*1e6+1.1567E-15*lr*1e6-3.068E-16))*nf+((-3.2841E-18*lr*lr*1e6*1e6+1.3358E-17*lr*1e6+1.7142E-17)*wr*wr*1e6*1e6+(5.3662E-17*lr*1e6*lr*1e6-2.4561E-16*lr*1e6-3.1695E-16)*wr*1e6+(-3.2421E-16*lr*lr*1e6*1e6+1.5991E-16*lr*1e6+3.211E-16)),1e-18)'
+Djdb_AREA_rf = '(nf/2*wr*(0.8-2*0.065))*1e-6'
+Djdb_PJ_rf   = '(1+1.7977e-7/wr)*nf*wr'
+Djsb_AREA_rf = '(wr*(0.8-0.065)*2+(nf/2-1)*wr*(0.8-2*0.065))*1e-6'
+Djsb_PJ_rf   = '(1+1.7977e-7/wr)*nf*wr'
+Rdc_n33_rf      = 'max((86.7923*exp(-0.1713*wr*1e6)),1e-3)'
+Rsc_n33_rf      =  'max((86.7923*exp(-0.1713*wr*1e6)),1e-3)'
+Rsub1_rf      = 'max(((0.0011*pwr(lr*1e6,0.0699)*log(wr*1e6))+(0.0064*pwr(lr*1e6,-0.1022)))*nf*nf+((-0.0197*log(lr*1e6)-0.0762)*wr*1e6+(0.2539*log(lr*1e6)-1.3244))*nf+((9.2323*lr*lr*1e6*1e6-16.353*lr*1e6+16.212)*wr*1e6+(103.21*lr*lr*1e6*1e6-183.88*lr*1e6+170.1)),1e-3)'
+Rsub2_rf      = 'max((0.0226*nf*nf-5.6376*nf+401.39),1e-3)'
+Rsub3_rf      = 'max((3062.5*pwr(nf,-0.8254)),1e-3)'
+Cgdo_n33_rf     = 'max((0+DCGDO_N33_RF),0)'
+Cgso_n33_rf     = 'max((0+DCGSO_N33_RF),0)'
+Cj_n33_rf    = 'max((0+dcj_n33_rf), 0)'
+Cjsw_n33_rf     = 'max((0+dcjsw_n33_rf), 0)'
*****************************************
Lgate       2 20 1p
Rgate       20 21 Rg_rf
Cgd_ext     20 11 Cgd_rf
Cgs_ext     20 31 Cgs_rf
Cds_ext     15 31 Cds_rf
Rds         11 15 1m
Ldrain      1 11 1p
Lsource     3 31 1p
*****************************************
Djdb  12 11
+ ndio33_rf
+ AREA  = Djdb_AREA_rf
+ PJ    = Djdb_PJ_rf 
***
Djsb  32 31
+ ndio33_rf
+ AREA  = Djsb_AREA_rf
+ PJ    = Djsb_PJ_rf
*****************************************
Rsub1      41  4  Rsub1_rf
Rsub2      41  12 Rsub2_rf
Rsub3      41  32 Rsub3_rf
*
* --------- ideal mos transistor ----------------------
MAIN 11 21 31 41 n33_rf L=lr W=wr m=nf AD = 0 AS = 0 PD = 0 PS = 0
* MOS Model
.MODEL n33_rf NMOS
+LEVEL = 49
*
* GENERAL PARAMETERS
*
+CALCACM  = 1
+LMIN     = 3.3E-7              LMAX     = 1.2E-6              WMIN     = 4.8E-7              
+WMAX     = 1.002E-5            TNOM     = 25.0                VERSION  = 3.24                 
+TOX      = '6.65E-09+DTOX_N33_RF' TOXM     = 6.65E-09            XJ       = 1.6000000E-07       
+NCH      = 4.3441000E+17       LLN      = 1.0625758           LWN      = 1.0101005           
+WLN      = 0.9810000           WWN      = 0.9060000           LINT     = 6.3891300E-08       
+LL       = -2.3305548E-15      LW       = -2.4634918E-15      LWL      = 2.6243002E-24       
+WINT     = 3.5850000E-08       WL       = -1.8902563E-15      WW       = -1.3000000E-14      
+WWL      = -1.3027796E-20      MOBMOD   = 1                   BINUNIT  = 2                   
+XL       = '1E-8+DXL_N33_RF'   XW       = '0.00+DXW_N33_RF'   DWG      = -3.9100000E-09                  
+DWB      = 3.2000000E-09       
* DIODE PARAMETERS
+ACM      = 12                  LDIF     = 6.50E-08            HDIF     = 2.05E-07            
+RSH      = 7.08                RD       = 0                   RS       = 0                   
+RSC      = 'Rsc_n33_rf'          RDC      =  'Rdc_n33_rf'                 
*
* THRESHOLD VOLTAGE PARAMETERS
*
+VTH0     = '0.695+DVTH_N33_RF'    LVTH0    = 4.0100000E-10       WVTH0    = 1.0200000E-08       
+PVTH0    = '8.0000000E-16+DPVTH0_N33_RF'       K1       = 0.8451000           LK1      = 5.8182560E-10       
+WK1      = -6.2456240E-09      PK1      = 1.9938927E-15       K2       = 4.4575000E-02       
+K3       = -3.8500000          DVT0     = 9.4991400           LDVT0    = 8.0839730E-09       
+DVT1     = 0.6300000           LDVT1    = 5.5000000E-08       DVT2     = -0.1450000          
+DVT0W    = 0.00                DVT1W    = 0.1057000           DVT2W    = 0.00                
+NLX      = 2.0274594E-07       LNLX     = -2.8608589E-14      W0       = 0.00                
+K3B      = 0.5669292           NGATE    = 2.6812141E+21                 
*
* MOBILITY PARAMETERS
*
+VSAT     = 8.5000000E+04       LVSAT    = -1.7300000E-03      PVSAT    = 1.2000000E-10       
+UA       = -8.6001130E-10      UB       = 2.3000001E-18       UC       = 1.3100000E-10       
+PUC      = 5.0000000E-25       RDSW     = 2.4208382E+02       PRWB     = -8.5000000E-02      
+PRWG     = 3.8000000E-02       WR       = 1.0000000           U0       = 3.5000000E-02       
+LU0      = 5.0000000E-10       A0       = 1.0200000           LA0      = -1.2000000E-07      
+KETA     = 0.00                LKETA    = -1.4000000E-08      WKETA    = -1.9999999E-09      
+PKETA    = 1.0000000E-15       A1       = 0.00                A2       = 0.9900000           
+AGS      = 0.1700000           B0       = 1.0000000E-08       B1       = 0.00                
*
* SUBTHRESHOLD CURRENT PARAMETERS
*
+VOFF     = -0.1200000          NFACTOR  = 1.1000000           LNFACTOR = 4.0000000E-08       
+PNFACTOR = -1.4000000E-14      CIT      = 1.0000000E-04       CDSC     = 5.0000000E-04       
+CDSCB    = 0.00                CDSCD    = 0.00                ETA0     = 4.0000000E-02       
+PETA0    = 3.0000001E-16       ETAB     = -0.1000000          DSUB     = 0.6000000           
*
* ROUT PARAMETERS
*
+PCLM     = 0.8000000           LPCLM    = 5.0000000E-08       PPCLM    = 8.0000000E-15       
+PDIBLC1  = 9.0000000E-02       PDIBLC2  = 1.6000000E-03       PPDIBLC2 = -7.0000000E-17      
+PDIBLCB  = 0.00                DROUT    = 0.5987002           PSCBE1   = 3.4000000E+08       
+LPSCBE1  = 13.0000000          PSCBE2   = 3.8000000E-06       PVAG     = 0.00                
+DELTA    = 1.0000000E-02       ALPHA0   = -4.4760000E-08      ALPHA1   = 0.8998877           
+BETA0    = 18.8771250          LBETA0   = -5.7118000E-07
*
* TEMPERATURE EFFECTS PARAMETERS
*
+KT1      = -0.3250000          PKT1     = -2.3708420E-15      KT2      = -3.6844640E-02      
+AT       = 2.2000000E+04       UTE      = -1.4100000          UA1      = 2.0599999E-09       
+WUA1     = -1.2600000E-16      PUA1     = -1.0000000E-24      UB1      = -2.5000000E-18      
+WUB1     = 1.1000000E-25       UC1      = -1.1000000E-10      LUC1     = 1.6999999E-17       
+KT1L     = -5.0000000E-09      PRT      = 40.0000000          
*
* CAPACITANCE PARAMETERS
*
+CJ       = 'Cj_n33_rf '                   MJ       = 0.321               PB       = 0.708               
+CJSW     = 'Cjsw_n33_rf'                   MJSW     = 0.447               PBSW     = 1                   
+CJSWG    = 0                   MJSWG    = 0.447               PBSWG    = 1                   
+TPB      = 0.00166             TPBSW    = 0.00162             TPBSWG   = 0.00162     
+TCJ      = 0.000897            TCJSW    = 0.000695            TCJSWG   = 0.000695
+JS       = 3.65E-07            JSW      = 3.0E-13             NJ       = 1.04                 
+XTI      = 3.9                 NQSMOD   = 0                   ELM      = 5 
+CGDO     = 'Cgdo_n33_rf'          CGSO     = 'Cgso_n33_rf'  CGBO = 0  TLEVC    = 1 
+CAPMOD   = 3                   XPART    = 1                   CF       = 0.00                  
+ACDE     = 0.45                MOIN     = 24                  NOFF     = 2.3177            
+DLC      = 6.50E-08            
*    
* NOISE PARAMETERS
*
+NOIMOD   = 2                   NOIA     = 1.5500E+20            NOIB     = 7.1866E+04    
+NOIC     = 1.4952E-13          EM       = 3.2163E+07            EF       = 9.9600E-01 
*
* Diode Model 
.MODEL ndio33_rf D
*
+LEVEL    = 3                   JS       = 3.65E-07            JSW      = 1E-15            
+N        = 1.0203              RS       = 8.84E-09            IK       = 1.33E+05            
+IKR      = 2.78E+05            BV       = 11.0                IBV      = 277.78              
+TRS      = 1.07E-03            EG       = 1.16                TREF     = 25.0                
+XTI      = 3.0                 CJ       = 0.000845            MJ       = 0.321               
+PB       = 0.708               CJSW     = 3.41E-10            MJSW     = 0.447               
+PHP      = 1                   CTA      = 0.000897            CTP      = 0.000695            
+TPB      = 0.00166             TPHP     = 0.00162             TLEV     = 1
+TLEVC    = 1                   AREA     = 3.60E-09            PJ       = 2.4E-04
+FC       = 0                   FCS      = 0  
.ends n33_ckt_rf
***************************
* 3.3V RF DNWMOS Subcircuit
***************************
* 11=drain, 2=gate, 31=source, 4=bulk
* lr=gate length, wr=finger width, nf=finger number, laddr=DNW diode add length, waddr=DNW diode add width
.subckt dnw33_ckt_rf 1 2 3 4 5 lr=l wr=w nf=finger laddr=ladd waddr=wadd
* scalable unit parameter
* euqivalent circuit saclable parameter
.param
+Rg_rf        = 'max((((337.44*lr*lr*1e6*1e6-636.15*lr*1e6+1247.8)*pwr(wr*1e6,(0.0345*lr*lr*1e6*1e6-0.0673*lr*1e6-0.8144)))*pwr(nf,(0.01549*lr*lr*1e6*1e6-0.02983*lr*1e6+0.10754)*log(wr*1e6)+(-0.01723*lr*lr*1e6*1e6+0.03465*lr*1e6-0.95262))),1e-3)'
+Cgd_rf       = 'max((((-1.019487e-18*lr*lr*1e6*1e6+2.093231E-18*lr*1e6-5.621744E-18)*wr*wr*1e6*1e6+(-7.0297E-17*lr*lr*1e6*1e6+1.4369E-16*lr*1e6+3.8644E-16)*wr*1e6+(9.4974E-18*lr*lr*1e6*1e6+3.9394E-17*lr*1e6+2.3454E-16))*nf+((-4.8156E-18*lr*lr*1e6*1e6+1.1596E-16*lr*1e6-2.1673E-17)*wr*wr*1e6*1e6+(4.816E-16*lr*lr*1e6*1e6-1.2046E-15*lr*1e6+8.1E-19)*wr*1e6+(-1.5056E-16*lr*lr*1e6*1e6+7.2245E-16*lr*1e6+2.1267E-16))),1e-18)'
+Cgs_rf       = 'max(((-1.7423e-17*lr*lr*1e6*1e6+3.3616E-17*lr*1e6+7.4972E-19)*wr*wr*1e6*1e6+(-8.3169E-17*lr*lr*1e6*1e6+2.8529E-16*lr*1e6+2.5325E-16)*wr*1e6+(-5.1487E-16*lr*lr*1e6*1e6+9.9831E-16*lr*1e6+3.2256E-16))*nf+((-2.5956E-17*lr*lr*1e6*1e6-2.5684E-17*lr*1e6+1.5362E-16)*wr*wr*1e6*1e6+(-3.6262E-15*lr*lr*1e6*1e6+6.3722E-15*lr*1e6-3.7861E-15)*wr*1e6+(8.4615E-15*lr*lr*1e6*1e6-1.4192E-14*lr*1e6+7.9308E-15)),1e-18)'
+Cds_rf       = 'max(((-8.3173e-17*lr*lr*1e6*1e6+1.4664E-16*lr*1e6-3.1474E-17)*wr*wr*1e6*1e6+(4.9488E-16*lr*lr*1e6*1e6-8.6038E-16*lr*1e6+4.8447E-16)*wr*1e6+(-6.5021E-16*lr*lr*1e6*1e6+1.1567E-15*lr*1e6-3.068E-16))*nf+((-3.2841E-18*lr*lr*1e6*1e6+1.3358E-17*lr*1e6+1.7142E-17)*wr*wr*1e6*1e6+(5.3662E-17*lr*1e6*lr*1e6-2.4561E-16*lr*1e6-3.1695E-16)*wr*1e6+(-3.2421E-16*lr*lr*1e6*1e6+1.5991E-16*lr*1e6+3.211E-16)),1e-18)'
+Djdb_AREA_rf = '(nf/2*wr*(0.8-2*0.065))*1e-6'
+Djdb_PJ_rf   = '(1+1.7977e-7/wr)*nf*wr'
+Djsb_AREA_rf = '(wr*(0.8-0.065)*2+(nf/2-1)*wr*(0.8-2*0.065))*1e-6'
+Djsb_PJ_rf   = '(1+1.7977e-7/wr)*nf*wr'
+Djbdn_AREA_rf= '(2*0.8*1e-6+lr*nf+0.8*1e-6*(nf-1)+2*laddr)*(wr+2*waddr)'
+Djbdn_PJ_rf  = '2*(2*0.8*1e-6+lr*nf+0.8*1e-6*(nf-1)+wr+2*(laddr+waddr))'
+Rdc_n33_rf      = 'max((86.7923*exp(-0.1713*wr*1e6)),1e-3)'
+Rsc_n33_rf      = 'max((86.7923*exp(-0.1713*wr*1e6)),1e-3)'
+Rsub1_rf      = 'max(((0.0011*pwr(lr*1e6,0.0699)*log(wr*1e6))+(0.0064*pwr(lr*1e6,-0.1022)))*nf*nf+((-0.0197*log(lr*1e6)-0.0762)*wr*1e6+(0.2539*log(lr*1e6)-1.3244))*nf+((9.2323*lr*lr*1e6*1e6-16.353*lr*1e6+16.212)*wr*1e6+(103.21*lr*lr*1e6*1e6-183.88*lr*1e6+170.1)),1e-3)'
+Rsub2_rf      = 'max((0.0226*nf*nf-5.6376*nf+401.39),1e-3)'
+Rsub3_rf      = 'max((3062.5*pwr(nf,-0.8254)),1e-3)'
+Cgdo_n33_rf     = 'max((0+DCGDO_N33_RF),0)'
+Cgso_n33_rf     = 'max((0+DCGSO_N33_RF),0)'
+Cj_n33_rf    = 'max((0+dcj_n33_rf), 0)'
+Cjsw_n33_rf     = 'max((0+dcjsw_n33_rf), 0)'
*****************************************
Lgate       2 20 1p
Rgate       20 21 Rg_rf
Cgd_ext     20 11 Cgd_rf
Cgs_ext     20 31 Cgs_rf
Cds_ext     15 31 Cds_rf
Rds         11 15 1m
Ldrain      1 11 1p
Lsource     3 31 1p
*****************************************
Djdb  12 11
+ ndio33_rf
+ AREA  = Djdb_AREA_rf
+ PJ    = Djdb_PJ_rf 
***
Djsb  32 31
+ ndio33_rf
+ AREA  = Djsb_AREA_rf
+ PJ    = Djsb_PJ_rf
***
Djbdn  4 5
+ diobpw_rf
+ AREA  = Djbdn_AREA_rf
+ PJ    = Djbdn_PJ_rf
*****************************************
Rsub1      41  4   Rsub1_rf
Rsub2      41  12  Rsub2_rf
Rsub3      41  32  Rsub3_rf
*
* --------- ideal mos transistor ----------------------
MAIN 11 21 31 41 dnw33_rf L=lr W=wr m=nf AD = 0 AS = 0 PD = 0 PS = 0
* MOS Model
.MODEL dnw33_rf NMOS
+LEVEL = 49
*
* GENERAL PARAMETERS
*
+CALCACM  = 1
+LMIN     = 3.3E-7              LMAX     = 1.2E-6              WMIN     = 4.8E-7              
+WMAX     = 1.002E-5            TNOM     = 25.0                VERSION  = 3.24                 
+TOX      = '6.65E-09+DTOX_N33_RF' TOXM     = 6.65E-09            XJ       = 1.6000000E-07       
+NCH      = 4.3441000E+17       LLN      = 1.0625758           LWN      = 1.0101005           
+WLN      = 0.9810000           WWN      = 0.9060000           LINT     = 6.3891300E-08       
+LL       = -2.3305548E-15      LW       = -2.4634918E-15      LWL      = 2.6243002E-24       
+WINT     = 3.5850000E-08       WL       = -1.8902563E-15      WW       = -1.3000000E-14      
+WWL      = -1.3027796E-20      MOBMOD   = 1                   BINUNIT  = 2                   
+XL       = '1E-8+DXL_N33_RF'   XW       = '0.00+DXW_N33_RF'   DWG      = -3.9100000E-09                  
+DWB      = 3.2000000E-09       
* DIODE PARAMETERS
+ACM      = 12                  LDIF     = 6.50E-08            HDIF     = 2.05E-07            
+RSH      = 7.08                RD       = 0                   RS       = 0                   
+RSC      = 'Rdc_n33_rf'           RDC      = 'Rdc_n33_rf'                 
*
* THRESHOLD VOLTAGE PARAMETERS
*
+VTH0     = '0.695+DVTH_N33_RF'    LVTH0    = 4.0100000E-10       WVTH0    = 1.0200000E-08       
+PVTH0    = '8.0000000E-16+DPVTH0_N33_RF'       K1       = 0.8451000           LK1      = 5.8182560E-10       
+WK1      = -6.2456240E-09      PK1      = 1.9938927E-15       K2       = 4.4575000E-02       
+K3       = -3.8500000          DVT0     = 9.4991400           LDVT0    = 8.0839730E-09       
+DVT1     = 0.6300000           LDVT1    = 5.5000000E-08       DVT2     = -0.1450000          
+DVT0W    = 0.00                DVT1W    = 0.1057000           DVT2W    = 0.00                
+NLX      = 2.0274594E-07       LNLX     = -2.8608589E-14      W0       = 0.00                
+K3B      = 0.5669292           NGATE    = 2.6812141E+21                 
*
* MOBILITY PARAMETERS
*
+VSAT     = 8.5000000E+04       LVSAT    = -1.7300000E-03      PVSAT    = 1.2000000E-10       
+UA       = -8.6001130E-10      UB       = 2.3000001E-18       UC       = 1.3100000E-10       
+PUC      = 5.0000000E-25       RDSW     = 2.4208382E+02       PRWB     = -8.5000000E-02      
+PRWG     = 3.8000000E-02       WR       = 1.0000000           U0       = 3.5000000E-02       
+LU0      = 5.0000000E-10       A0       = 1.0200000           LA0      = -1.2000000E-07      
+KETA     = 0.00                LKETA    = -1.4000000E-08      WKETA    = -1.9999999E-09      
+PKETA    = 1.0000000E-15       A1       = 0.00                A2       = 0.9900000           
+AGS      = 0.1700000           B0       = 1.0000000E-08       B1       = 0.00                
*
* SUBTHRESHOLD CURRENT PARAMETERS
*
+VOFF     = -0.1200000          NFACTOR  = 1.1000000           LNFACTOR = 4.0000000E-08       
+PNFACTOR = -1.4000000E-14      CIT      = 1.0000000E-04       CDSC     = 5.0000000E-04       
+CDSCB    = 0.00                CDSCD    = 0.00                ETA0     = 4.0000000E-02       
+PETA0    = 3.0000001E-16       ETAB     = -0.1000000          DSUB     = 0.6000000           
*
* ROUT PARAMETERS
*
+PCLM     = 0.8000000           LPCLM    = 5.0000000E-08       PPCLM    = 8.0000000E-15       
+PDIBLC1  = 9.0000000E-02       PDIBLC2  = 1.6000000E-03       PPDIBLC2 = -7.0000000E-17      
+PDIBLCB  = 0.00                DROUT    = 0.5987002           PSCBE1   = 3.4000000E+08       
+LPSCBE1  = 13.0000000          PSCBE2   = 3.8000000E-06       PVAG     = 0.00                
+DELTA    = 1.0000000E-02       ALPHA0   = -4.4760000E-08      ALPHA1   = 0.8998877           
+BETA0    = 18.8771250          LBETA0   = -5.7118000E-07
*
* TEMPERATURE EFFECTS PARAMETERS
*
+KT1      = -0.3250000          PKT1     = -2.3708420E-15      KT2      = -3.6844640E-02      
+AT       = 2.2000000E+04       UTE      = -1.4100000          UA1      = 2.0599999E-09       
+WUA1     = -1.2600000E-16      PUA1     = -1.0000000E-24      UB1      = -2.5000000E-18      
+WUB1     = 1.1000000E-25       UC1      = -1.1000000E-10      LUC1     = 1.6999999E-17       
+KT1L     = -5.0000000E-09      PRT      = 40.0000000          
*
* CAPACITANCE PARAMETERS
*
+CJ       = 'Cj_n33_rf'                  MJ       = 0.321               PB       = 0.708               
+CJSW     = 'Cjsw_n33_rf'                   MJSW     = 0.447               PBSW     = 1                   
+CJSWG    = 0                   MJSWG    = 0.447               PBSWG    = 1                   
+TPB      = 0.00166             TPBSW    = 0.00162             TPBSWG   = 0.00162     
+TCJ      = 0.000897            TCJSW    = 0.000695            TCJSWG   = 0.000695
+JS       = 3.65E-07            JSW      = 3.0E-13             NJ       = 1.04                 
+XTI      = 3.9                 NQSMOD   = 0                   ELM      = 5 
+CGDO     = 'Cgdo_n33_rf'          CGSO     = 'Cgso_n33_rf'   CGBO = 0       TLEVC    = 1 
+CAPMOD   = 3                   XPART    = 1                   CF       = 0.00                  
+ACDE     = 0.45                MOIN     = 24                  NOFF     = 2.3177            
+DLC      = 6.50E-08            
*    
* NOISE PARAMETERS
*
+NOIMOD   = 2                   NOIA     = 1.5500E+20            NOIB     = 7.1866E+04    
+NOIC     = 1.4952E-13          EM       = 3.2163E+07            EF       = 9.9600E-01 
*
* Diode Model 
.MODEL ndio33_rf D
*
+LEVEL    = 3                   JS       = 3.65E-07            JSW      = 1E-15            
+N        = 1.0203              RS       = 8.84E-09            IK       = 1.33E+05            
+IKR      = 2.78E+05            BV       = 11.0                IBV      = 277.78              
+TRS      = 1.07E-03            EG       = 1.16                TREF     = 25.0                
+XTI      = 3.0                 CJ       = 0.000845            MJ       = 0.321               
+PB       = 0.708               CJSW     = 3.41E-10            MJSW     = 0.447               
+PHP      = 1                   CTA      = 0.000897            CTP      = 0.000695            
+TPB      = 0.00166             TPHP     = 0.00162             TLEV     = 1
+TLEVC    = 1                   AREA     = 3.60E-09            PJ       = 2.4E-04
+FC       = 0                   FCS      = 0 
* Diode Model  
.model diobpw_rf D
*    
+LEVEL    = 3                   JS       = 1.50E-07            JSW      = 1.00E-15            
+N        = 1.0213              RS       = 2.51E-08            IK       = 2.40E+05            
+IKR      = 1.04E+05            BV       = 15.0                IBV      = 1.04E+02                
+TRS      = 1.77E-03            CTA      = 0.0012              CTP      = 0.00107                
+EG       = 1.16                TREF     = 25.0                TPB      = 0.0019               
+TPHP     = 0.00193             XTI      = 3.0                 CJ       = 0.000536            
+MJ       = 0.343               PB       = 0.693               CJSW     = 3.22E-10            
+MJSW     = 0.361               PHP      = 0.715               TLEV     = 1
+TLEVC    = 1      		AREA     = 9.6E-9              PJ       = 4E-4  
+FC       = 0                   FCS      = 0
.ends dnw33_ckt_rf
*************************
* 3.3V RF PMOS Subcircuit
*************************
* 11=drain, 2=gate, 31=source, 4=bulk
* lr=gate length, wr=finger width, nf=finger number
.subckt p33_ckt_rf 1 2 3 4 lr=l wr=w nf=finger
* scalable unit parameter
* euqivalent circuit saclable parameter
.param
+Rg_rf        = 'max(((-0.1307*pwr(lr*1e6,2)-0.1679*lr*1e6+0.3067)*pwr(wr*1e6,2)+(-1.5879*pwr(lr*1e6,2)+6.3308*lr*1e6-4.3942)*wr*1e6+(0.1019*pwr(lr*1e6,2)-17.347*lr*1e6+14.299))+((-110.36*pwr(lr*1e6,2)+173.06*lr*1e6-51.853)*pwr(wr*1e6,2)+(1223.8*pwr(lr*1e6,2)-1968.5*lr*1e6+557.24)*wr*1e6+(-988.57*pwr(lr*1e6,2)+2030.6*lr*1e6-114))/NF,1e-3)'
+Cgd_rf       = 'max((((0.0069*pwr(lr*1e6,2)-0.006*lr*1e6+0.0012)*pwr(wr*1e6,2)+(-0.05*pwr(lr*1e6,2)+0.0436*lr*1e6-0.0084)*wr*1e6+(0.0294*pwr(lr*1e6,2)-0.0285*lr*1e6+0.006))*Pwr(nf,2)+((-0.1241*pwr(lr*1e6,2)+0.1438*lr*1e6-0.0334)*pwr(wr*1e6,2)+(0.9454*pwr(lr*1e6,2)-1.0343*lr*1e6+0.5294)*wr*1e6+(-1.2623*pwr(lr*1e6,2)+1.5818*lr*1e6-0.085))*NF+((0.7611*pwr(lr*1e6,2)-1.0199*lr*1e6+0.2764)*pwr(wr*1e6,2)+(-7.3404*pwr(lr*1e6,2)+9.8018*lr*1e6-2.568)*wr*1e6+(10.408*pwr(lr*1e6,2)-14.261*lr*1e6+4.2573)))*1e-15,1e-18)'
+Cgs_rf       = 'max((((-0.0556*pwr(lr*1e6,2)+0.072*lr*1e6-0.0164)*pwr(wr*1e6,2)+(0.3886*pwr(lr*1e6,2)-0.5059*lr*1e6+0.1173)*wr*1e6+(-0.563*pwr(lr*1e6,2)+0.7329*lr*1e6-0.1699))*Pwr(nf,2)+((0.3657*pwr(lr*1e6,2)-0.4886*lr*1e6+0.1229)*pwr(wr*1e6,2)+(-3.0209*pwr(lr*1e6,2)+3.4127*lr*1e6-0.6043)*wr*1e6+(6.3133*pwr(lr*1e6,2)-8.2461*lr*1e6+2.374))*NF+((-0.777*pwr(lr*1e6,2)+1.1371*lr*1e6-0.3601)*pwr(wr*1e6,2)+(2.2591*pwr(lr*1e6,2)-7.4763*lr*1e6+3.6663)*wr*1e6+(-6.6803*pwr(lr*1e6,2)+14.463*lr*1e6-3.2627)))*1e-15,1e-18)'
+Cds_rf       = 'max((((-0.0344*pwr(lr*1e6,2)+0.0349*lr*1e6-0.0075)*pwr(wr*1e6,2)+(0.3513*pwr(lr*1e6,2)-0.3435*lr*1e6+0.0732)*wr*1e6+(-0.5587*pwr(lr*1e6,2)+0.541*lr*1e6-0.115))*Pwr(nf,2)+((0.469*pwr(lr*1e6,2)-0.4217*lr*1e6+0.0652)*pwr(wr*1e6,2)+(-5.422*pwr(lr*1e6,2)+4.6966*lr*1e6-0.2819)*wr*1e6+(8.8347*pwr(lr*1e6,2)-8.0843*lr*1e6+1.5796))*NF+((-0.708*pwr(lr*1e6,2)+0.2244*lr*1e6+0.1665)*pwr(wr*1e6,2)+(9.9669*pwr(lr*1e6,2)-5.1155*lr*1e6-0.9422)*wr*1e6+(-16.183*pwr(lr*1e6,2)+9.5447*lr*1e6+1.0176)))*1e-15,1e-18)'
+Djdb_AREA_rf = '(nf/2*wr*1e6*(0.8-2*0.065))*1e-12'
+Djdb_PJ_rf   = '(0.99997+1.8823e-7/wr*1e6)*nf*wr'
+Djsb_AREA_rf = '(wr*1e6*(0.8-0.065)*2+(nf/2-1)*wr*1e6*(0.8-2*0.065))*1e-12'
+Djsb_PJ_rf   = '(0.99997+1.8823e-7/wr*1e6)*nf*wr'
+Rdc_p33      = 'max((300/(wr*1e6)), 1e-3)'
+Rsc_p33      = 'max((300/(wr*1e6)), 1e-3)'
+Cgdo_p33     = 'max((0+DCGDO_P33_RF),0)'
+Cgso_p33     = 'max((0+DCGSO_P33_RF),0)'
+Rds_rf       = 'max(((375.75*pwr(lr*1e6,2)-603.31*lr*1e6+131.78)*pwr(wr*1e6,2)+(-4158.8*pwr(lr*1e6,2)+6647.4*lr*1e6-1413.4)*wr*1e6+(5776.5*pwr(lr*1e6,2)-7973.7*lr*1e6+1834.2))*pwr(nf,(-0.085*pwr(lr*1e6,2)+0.1295*lr*1e6-0.0224)*pwr(wr*1e6,2)+(0.7499*pwr(lr*1e6,2)-1.2094*lr*1e6+0.1621)*wr*1e6+(-0.859*pwr(lr*1e6,2)+1.1497*lr*1e6-0.4753)), 1e-3)'
+Rsub2_rf     = 'max(((942147*pwr(lr*1e6,2)-1000000*lr*1e6+466678)*pwr(wr*1e6,2)+(-2000000*pwr(lr*1e6,2)+4000000*lr*1e6-1000000)*wr*1e6+(1000000*pwr(lr*1e6,2)-2000000*lr*1e6+873325))*pwr(nf,(-0.2537*pwr(lr*1e6,2)+0.354*lr*1e6-0.0821)*pwr(wr*1e6,2)+(1.3061*pwr(lr*1e6,2)-1.8324*lr*1e6+0.1598)*wr*1e6+(-1.0001*pwr(lr*1e6,2)+1.4236*lr*1e6-0.2592)), 1e-3)'
+Rsub3_rf     = 'max(((942147*pwr(lr*1e6,2)-1000000*lr*1e6+466678)*pwr(wr*1e6,2)+(-2000000*pwr(lr*1e6,2)+4000000*lr*1e6-1000000)*wr*1e6+(1000000*pwr(lr*1e6,2)-2000000*lr*1e6+873325))*pwr(nf,(-0.2537*pwr(lr*1e6,2)+0.354*lr*1e6-0.0821)*pwr(wr*1e6,2)+(1.3061*pwr(lr*1e6,2)-1.8324*lr*1e6+0.1598)*wr*1e6+(-1.0001*pwr(lr*1e6,2)+1.4236*lr*1e6-0.2592)), 1e-3)'
+Cj_p33       = 'max((0+dcj_p33_rf), 0)'
+Cjsw_p33     = 'max((0+dcjsw_p33_rf), 0)'
*****************************************
Lgate       2 20  1p
Rgate       20 21 Rg_rf
Cgd_ext     20 11 Cgd_rf
Cgs_ext     20 31 Cgs_rf
Cds_ext     15 31 Cds_rf
Rds         11 15 Rds_rf
Ldrain       1 11 1p
Lsource      3 31 1p
*****************************************
Djdb  11 12
+ pdio33_rf
+ AREA  = Djdb_AREA_rf
+ PJ    = Djdb_PJ_rf 
***
Djsb  31 32
+ pdio33_rf
+ AREA  = Djsb_AREA_rf
+ PJ    = Djsb_PJ_rf
*****************************************
Rsub1      41  4  3
Rsub2      41  12 Rsub2_rf
Rsub3      41  32 Rsub3_rf
*
* --------- ideal mos transistor ----------------------
MAIN 11 21 31 41 p33_rf L=lr W=wr m=nf AD = 0 AS = 0 PD = 0 PS = 0
* MOS Model
.MODEL p33_rf PMOS
+LEVEL = 49
*
* GENERAL PARAMETERS
*
+CALCACM  = 1
+LMIN     = 2.8E-7              LMAX     = 1.2E-6              WMIN     = 4.8E-7              
+WMAX     = 1.002E-5            TNOM     = 25.0                VERSION  = 3.24                 
+TOX      = '6.62E-09+DTOX_P33_RF' TOXM     = 6.62E-09            XJ       = 1.7000001E-07       
+NCH      = 5.4852000E+17       LLN      = 1.0471729           LWN      = 0.9530895           
+WLN      = 1.0257638           WWN      = 0.9617700           LINT     = 3.5000000E-08       
+LL       = 5.5000000E-15       LW       = -4.7160380E-14      LWL      = 7.0054450E-22       
+WINT     = 1.3000000E-08       WL       = -3.1491245E-14      WW       = 2.3000000E-15       
+WWL      = -2.4167156E-22      MOBMOD   = 1                   BINUNIT  = 2                   
+XL       = '-1.70E-08+DXL_P33_RF' XW       = '0.00+DXW_P33_RF'      DWG      = 0.00                   
+DWB      = 8.6000000E-09                                 
* DIODE PARAMETERS
+ACM      = 12                  LDIF     = 6.50E-08            HDIF     = 2.05E-07            
+RSH      = 9.8                 RD       = 0                   RS       = 0                   
+RSC      = 'Rsc_p33'           RDC      = 'Rdc_p33'                   
*
* THRESHOLD VOLTAGE PARAMETERS
*
+VTH0     = '-0.672+DVTH_P33_RF'   WVTH0    = 4.0000000E-09       PVTH0    = '6.0000000E-15+DPVTH0_P33_RF'       
+K1       = 0.9145741           PK1      = -1.7000000E-14      K2       = 4.1276220E-02       
+K3       = 0.1293833           DVT0     = 1.8000000           DVT1     = 0.7100000           
+DVT2     = -7.0000000E-02      DVT0W    = 0.00                DVT1W    = 0.00                
+DVT2W    = 0.00                NLX      = 1.2000000E-08       W0       = 1.0021131E-09       
+K3B      = 0.4000000           NGATE    = 1.1600000E+20               
*
* MOBILITY PARAMETERS
*
+VSAT     = 8.5500000E+04       PVSAT    = -5.8000000E-09      UA       = 3.1500000E-10       
+LUA      = 1.5000001E-17       WUA      = -1.6763224E-16      PUA      = -1.1000000E-23      
+UB       = 1.0444180E-18       LUB      = -7.0000000E-27      UC       = -3.5000000E-11      
+LUC      = 4.0000000E-18       PUC      = 5.0000000E-24       RDSW     = 9.5000000E+02       
+PRWB     = 0.00                PRWG     = 6.3755660E-03       WR       = 1.0000000           
+U0       = 9.2500000E-03       LU0      = -4.1500680E-10      WU0      = -1.7001526E-12      
+PU0      = -3.7999640E-16      A0       = 0.8500000           KETA     = 1.5000000E-02       
+LKETA    = -1.0000000E-08      WKETA    = 1.0000000E-09       PKETA    = -6.0000000E-15      
+A1       = 0.00                A2       = 0.9900000           AGS      = 4.0000000E-02       
+B0       = 4.6000000E-08       B1       = 0.00                
*
* SUBTHRESHOLD CURRENT PARAMETERS
*
+VOFF     = -0.1000000          LVOFF    = 1.8000000E-09       PVOFF    = -2.9999999E-15      
+NFACTOR  = 1.1000000           PNFACTOR = -4.0000000E-14      CIT      = 1.9999999E-04       
+CDSC     = 4.5263850E-05       CDSCB    = 0.00                CDSCD    = 0.00                
+ETA0     = 5.0000000E-03       PETA0    = 7.0000000E-15       ETAB     = -1.5000000E-02      
+PETAB    = -2.0000000E-15      DSUB     = 0.5800000           
*
* ROUT PARAMETERS
*
+PCLM     = 0.6000000           PPCLM    = 1.3000000E-13       PDIBLC1  = 6.0000000E-03       
+PDIBLC2  = 2.5000001E-04       WPDIBLC2 = 8.0000000E-11       PDIBLCB  = 0.00                
+DROUT    = 0.5600000           PSCBE1   = 3.3000000E+08       PPSCBE1  = -7.0000000E-06      
+PSCBE2   = 2.0000000E-07       PVAG     = 0.00                DELTA    = 8.0000000E-03       
+PDELTA   = 4.0000000E-16       ALPHA0   = 1.3410400E-06       ALPHA1   = 5.6136910E-02       
+BETA0    = 27.5998000          
*
* TEMPERATURE EFFECTS PARAMETERS
*
+KT1      = -0.3840900          WKT1     = -9.4333370E-10      PKT1     = 4.9999980E-15       
+KT2      = -4.1563480E-02      AT       = -2.0000000E+03      PAT      = -7.5000000E-09      
+UTE      = -1.3236057          UA1      = 3.0000002E-10       WUA1     = 8.0000000E-18       
+PUA1     = 1.0000000E-23       UB1      = -2.0704662E-18      WUB1     = 1.4000000E-25       
+UC1      = -5.0000000E-11      KT1L     = -6.0000000E-09      PRT      = 1.3000000E+02
*
* CAPACITANCE PARAMETERS
*
+CJ       = 'Cj_p33'               MJ       = 0.401                PB       = 0.807
+CJSW     = 'Cjsw_p33'             MJSW     = 0.45                 PBSW     = 1
+CJSWG    = 0                      MJSWG    = 0.45                 PBSWG    = 1
+TPB      = 0.00157                TPBSW    = 0.00137              TPBSWG   = 0.00137
+TCJ      = 0.000883               TCJSW    = 0.000709             TCJSWG   = 0.000709
+JS       = 1.68E-07               JSW      = 4.0E-13              NJ       = 1.07
+XTI      = 3.0                    NQSMOD   = 0                    ELM      = 5
+CGDO     = 'Cgdo_p33'             CGSO     = 'Cgso_p33'           TLEVC    = 1
+CAPMOD   = 3                      XPART    = 1                    CF       = 0.00
+ACDE     = 0.55                   MOIN     = 15                   NOFF     = 0.565
+DLC      = 7.0E-09                DWC      = 6.0E-8               CGBO=0
*
* NOISE PARAMETERS
*
+NOIMOD   = 2                   NOIA     = 3.5911E+19            NOIB     = 3.0215E+03    
+NOIC     = 6.7064E-12          EM       = 4.2400E+07            EF       = 1.0829E+00 
*
.MODEL pdio33_rf D
+LEVEL    = 3                   JS       = 1.68E-07            JSW      = 1E-15            
+N        = 1.0143              RS       = 0                   IK       = 4.07E+05            
+IKR      = 2.78E+05            BV       = 11.0                IBV      = 277.78              
+TRS      = 1.24E-03            EG       = 1.16                TREF     = 25.0                
+XTI      = 3.0                 CJ       = 0.00101             MJ       = 0.401               
+PB       = 0.807               CJSW     = 8.96E-11            MJSW     = 0.45                
+PHP      = 1                   CTA      = 0.000883            CTP      = 0.000709            
+TPB      = 0.00157             TPHP     = 0.00137             TLEV     = 1
+TLEVC    = 1                   FC       = 0                   FCS      = 0 
.ends p33_ckt_rf

